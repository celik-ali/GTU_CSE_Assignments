module temp_gen(output [31:0] temp, input [31:0] orig);// For copying a number to prevent permanent changes.
	
	and temp1  (temp[0], 1, orig[0]);
	and temp2  (temp[1], 1, orig[1]);
	and temp3  (temp[2], 1, orig[2]);
	and temp4  (temp[3], 1, orig[3]);
	and temp5  (temp[4], 1, orig[4]);
	and temp6  (temp[5], 1, orig[5]);
	and temp7  (temp[6], 1, orig[6]);
	and temp8  (temp[7], 1, orig[7]);
	and temp9  (temp[8], 1, orig[8]);
	and temp10 (temp[9], 1, orig[9]);
	and temp11 (temp[10], 1, orig[10]);
	and temp12 (temp[11], 1, orig[11]);
	and temp13 (temp[12], 1, orig[12]);
	and temp14 (temp[13], 1, orig[13]);
	and temp15 (temp[14], 1, orig[14]);
	and temp16 (temp[15], 1, orig[15]);
	and temp17 (temp[16], 1, orig[16]);
	and temp18 (temp[17], 1, orig[17]);
	and temp19 (temp[18], 1, orig[18]);
	and temp20 (temp[19], 1, orig[19]);
	and temp21 (temp[20], 1, orig[20]);
	and temp22 (temp[21], 1, orig[21]);
	and temp23 (temp[22], 1, orig[22]);
	and temp24 (temp[23], 1, orig[23]);
	and temp25 (temp[24], 1, orig[24]);
	and temp26 (temp[25], 1, orig[25]);
	and temp27 (temp[26], 1, orig[26]);
	and temp28 (temp[27], 1, orig[27]);
	and temp29 (temp[28], 1, orig[28]);
	and temp30 (temp[29], 1, orig[29]);
	and temp31 (temp[30], 1, orig[30]);
	and temp32 (temp[31], 1, orig[31]);

endmodule
