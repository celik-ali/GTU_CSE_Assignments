module memory_block(output reg [31:0] read_data, input byteOperations, input [17:0] address, input[31:0] write_data, input memRead, memWrite);
//Couldn't implement because I have started late.
endmodule
