module move(output[31:0] res, input [31:0] rs, rt);


endmodule

